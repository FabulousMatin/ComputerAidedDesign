module NOT (
    input  A,
    output out
);

  _ACT_C1 _NOT (
      1,
      1,
      1,
      0,
      0,
      0,
      A,
      0,
      out
  );

endmodule
