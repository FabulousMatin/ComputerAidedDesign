module AND3 (
    input A, B, C,

    output out
);

    _ACT_C1 and3(0, 0, 0, 0, C, B, A, 0, out);

endmodule